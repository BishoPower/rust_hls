// Generated for AMD Alveo U50 - PIPELINED VERSION (CLEAN)
// Pipeline: 3-stage complex logic implementation
// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

module hft_zero_plus #(
    parameter integer DATA_WIDTH = 32,
    parameter integer ADDR_WIDTH = 16
) (
    // Clock and Reset
    input  wire                    ap_clk,
    input  wire                    ap_rst_n,
    
    // Control signals (HLS-style)
    input  wire                    ap_start,
    output reg                     ap_done,
    output wire                    ap_idle,
    output wire                    ap_ready,
    
    // Data inputs
    input  wire [DATA_WIDTH-1:0]  best_bid_price,
    input  wire [DATA_WIDTH-1:0]  best_ask_price,
    input  wire [DATA_WIDTH-1:0]  best_bid_qty,
    input  wire [DATA_WIDTH-1:0]  best_ask_qty,
    input  wire [DATA_WIDTH-1:0]  bid_queue_strong,
    input  wire [DATA_WIDTH-1:0]  ask_queue_strong,
    input  wire [DATA_WIDTH-1:0]  current_position,
    input  wire [DATA_WIDTH-1:0]  last_fill_price,
    input  wire [DATA_WIDTH-1:0]  last_fill_side,
    
    // Data outputs
    output wire [DATA_WIDTH-1:0]  action,
    output wire [DATA_WIDTH-1:0]  price,
    output wire [DATA_WIDTH-1:0]  quantity
);

    // Complex computation pipeline
    // Intermediate computation wires
    wire [DATA_WIDTH-1:0] node_9;
    wire [DATA_WIDTH-1:0] node_11;
    wire [DATA_WIDTH-1:0] node_12;
    wire [DATA_WIDTH-1:0] node_14;
    wire [DATA_WIDTH-1:0] node_16;
    wire [DATA_WIDTH-1:0] node_17;
    wire [DATA_WIDTH-1:0] node_18;
    wire [DATA_WIDTH-1:0] node_19;
    wire [DATA_WIDTH-1:0] node_20;
    wire [DATA_WIDTH-1:0] node_21;
    wire [DATA_WIDTH-1:0] node_22;
    wire [DATA_WIDTH-1:0] node_26;
    wire [DATA_WIDTH-1:0] node_27;
    wire [DATA_WIDTH-1:0] node_28;
    wire [DATA_WIDTH-1:0] node_29;
    wire [DATA_WIDTH-1:0] node_32;
    wire [DATA_WIDTH-1:0] node_33;
    wire [DATA_WIDTH-1:0] node_37;
    wire [DATA_WIDTH-1:0] node_38;
    wire [DATA_WIDTH-1:0] node_39;
    wire [DATA_WIDTH-1:0] node_40;
    wire [DATA_WIDTH-1:0] node_41;
    wire [DATA_WIDTH-1:0] node_42;
    wire [DATA_WIDTH-1:0] node_43;
    wire [DATA_WIDTH-1:0] node_44;
    wire [DATA_WIDTH-1:0] node_45;
    wire [DATA_WIDTH-1:0] node_46;
    wire [DATA_WIDTH-1:0] node_47;
    wire [DATA_WIDTH-1:0] node_48;
    wire [DATA_WIDTH-1:0] node_49;
    wire [DATA_WIDTH-1:0] node_50;
    wire [DATA_WIDTH-1:0] node_51;
    wire [DATA_WIDTH-1:0] node_52;
    wire [DATA_WIDTH-1:0] node_53;
    wire [DATA_WIDTH-1:0] node_54;
    wire [DATA_WIDTH-1:0] node_55;
    wire [DATA_WIDTH-1:0] node_56;
    wire [DATA_WIDTH-1:0] node_57;
    wire [DATA_WIDTH-1:0] node_58;
    wire [DATA_WIDTH-1:0] node_59;
    wire [DATA_WIDTH-1:0] node_60;
    wire [DATA_WIDTH-1:0] node_61;
    wire [DATA_WIDTH-1:0] node_62;
    wire [DATA_WIDTH-1:0] node_63;
    wire [DATA_WIDTH-1:0] node_64;
    wire [DATA_WIDTH-1:0] node_65;
    wire [DATA_WIDTH-1:0] node_66;
    wire [DATA_WIDTH-1:0] node_67;
    wire [DATA_WIDTH-1:0] node_68;
    wire [DATA_WIDTH-1:0] node_69;
    wire [DATA_WIDTH-1:0] node_70;
    wire [DATA_WIDTH-1:0] node_71;
    wire [DATA_WIDTH-1:0] node_72;
    wire [DATA_WIDTH-1:0] node_73;
    wire [DATA_WIDTH-1:0] node_74;
    wire [DATA_WIDTH-1:0] node_75;
    wire [DATA_WIDTH-1:0] node_76;
    wire [DATA_WIDTH-1:0] node_77;
    wire [DATA_WIDTH-1:0] node_78;
    wire [DATA_WIDTH-1:0] node_79;
    wire [DATA_WIDTH-1:0] node_80;
    wire [DATA_WIDTH-1:0] node_81;
    wire [DATA_WIDTH-1:0] node_82;
    wire [DATA_WIDTH-1:0] node_83;
    wire [DATA_WIDTH-1:0] node_84;
    wire [DATA_WIDTH-1:0] node_85;
    wire [DATA_WIDTH-1:0] node_86;
    wire [DATA_WIDTH-1:0] node_87;
    wire [DATA_WIDTH-1:0] node_88;
    wire [DATA_WIDTH-1:0] node_89;
    wire [DATA_WIDTH-1:0] node_90;
    wire [DATA_WIDTH-1:0] node_91;
    wire [DATA_WIDTH-1:0] node_92;
    wire [DATA_WIDTH-1:0] node_93;
    wire [DATA_WIDTH-1:0] node_94;
    wire [DATA_WIDTH-1:0] node_95;
    wire [DATA_WIDTH-1:0] node_96;
    wire [DATA_WIDTH-1:0] node_97;
    wire [DATA_WIDTH-1:0] node_98;
    wire [DATA_WIDTH-1:0] node_99;
    wire [DATA_WIDTH-1:0] node_100;
    wire [DATA_WIDTH-1:0] node_101;
    wire [DATA_WIDTH-1:0] node_102;
    wire [DATA_WIDTH-1:0] node_103;
    wire [DATA_WIDTH-1:0] node_104;
    wire [DATA_WIDTH-1:0] node_105;
    wire [DATA_WIDTH-1:0] node_106;
    wire [DATA_WIDTH-1:0] node_107;
    wire [DATA_WIDTH-1:0] node_108;
    wire [DATA_WIDTH-1:0] node_109;
    wire [DATA_WIDTH-1:0] node_110;
    wire [DATA_WIDTH-1:0] node_111;
    wire [DATA_WIDTH-1:0] node_112;
    wire [DATA_WIDTH-1:0] node_113;
    wire [DATA_WIDTH-1:0] node_114;
    wire [DATA_WIDTH-1:0] node_115;
    wire [DATA_WIDTH-1:0] node_116;
    wire [DATA_WIDTH-1:0] node_117;
    wire [DATA_WIDTH-1:0] node_118;
    wire [DATA_WIDTH-1:0] node_119;
    wire [DATA_WIDTH-1:0] node_120;
    wire [DATA_WIDTH-1:0] node_121;
    wire [DATA_WIDTH-1:0] node_122;
    wire [DATA_WIDTH-1:0] node_123;
    wire [DATA_WIDTH-1:0] node_124;
    wire [DATA_WIDTH-1:0] node_125;
    wire [DATA_WIDTH-1:0] node_126;
    wire [DATA_WIDTH-1:0] node_127;
    wire [DATA_WIDTH-1:0] node_128;
    wire [DATA_WIDTH-1:0] node_129;
    wire [DATA_WIDTH-1:0] node_130;
    wire [DATA_WIDTH-1:0] node_131;
    wire [DATA_WIDTH-1:0] node_132;
    wire [DATA_WIDTH-1:0] node_133;
    wire [DATA_WIDTH-1:0] node_134;
    wire [DATA_WIDTH-1:0] node_135;
    wire [DATA_WIDTH-1:0] node_136;
    wire [DATA_WIDTH-1:0] node_137;
    wire [DATA_WIDTH-1:0] node_138;
    wire [DATA_WIDTH-1:0] node_139;
    wire [DATA_WIDTH-1:0] node_140;
    wire [DATA_WIDTH-1:0] node_141;
    wire [DATA_WIDTH-1:0] node_142;
    wire [DATA_WIDTH-1:0] node_143;
    wire [DATA_WIDTH-1:0] node_144;
    wire [DATA_WIDTH-1:0] node_145;
    wire [DATA_WIDTH-1:0] node_146;
    wire [DATA_WIDTH-1:0] node_147;
    wire [DATA_WIDTH-1:0] node_148;
    wire [DATA_WIDTH-1:0] node_149;
    wire [DATA_WIDTH-1:0] node_150;
    wire [DATA_WIDTH-1:0] node_151;
    wire [DATA_WIDTH-1:0] node_152;
    wire [DATA_WIDTH-1:0] node_153;
    wire [DATA_WIDTH-1:0] node_154;
    wire [DATA_WIDTH-1:0] node_155;
    wire [DATA_WIDTH-1:0] node_156;
    wire [DATA_WIDTH-1:0] node_157;
    wire [DATA_WIDTH-1:0] node_158;
    wire [DATA_WIDTH-1:0] node_159;
    wire [DATA_WIDTH-1:0] node_160;
    wire [DATA_WIDTH-1:0] node_161;
    wire [DATA_WIDTH-1:0] node_162;
    wire [DATA_WIDTH-1:0] node_163;
    wire [DATA_WIDTH-1:0] node_164;
    wire [DATA_WIDTH-1:0] node_165;
    wire [DATA_WIDTH-1:0] node_166;
    wire [DATA_WIDTH-1:0] node_167;
    wire [DATA_WIDTH-1:0] node_168;
    wire [DATA_WIDTH-1:0] node_169;
    wire [DATA_WIDTH-1:0] node_170;
    wire [DATA_WIDTH-1:0] node_171;
    wire [DATA_WIDTH-1:0] node_172;
    wire [DATA_WIDTH-1:0] node_173;
    wire [DATA_WIDTH-1:0] node_174;
    wire [DATA_WIDTH-1:0] node_175;
    wire [DATA_WIDTH-1:0] node_176;
    wire [DATA_WIDTH-1:0] node_177;
    wire [DATA_WIDTH-1:0] node_178;
    wire [DATA_WIDTH-1:0] node_179;
    wire [DATA_WIDTH-1:0] node_180;
    wire [DATA_WIDTH-1:0] node_181;
    wire [DATA_WIDTH-1:0] node_182;
    wire [DATA_WIDTH-1:0] node_183;
    wire [DATA_WIDTH-1:0] node_184;
    wire [DATA_WIDTH-1:0] node_185;
    wire [DATA_WIDTH-1:0] node_186;
    wire [DATA_WIDTH-1:0] node_187;
    wire [DATA_WIDTH-1:0] node_188;
    wire [DATA_WIDTH-1:0] node_189;
    wire [DATA_WIDTH-1:0] node_190;
    wire [DATA_WIDTH-1:0] node_191;
    wire [DATA_WIDTH-1:0] node_192;
    wire [DATA_WIDTH-1:0] node_193;
    wire [DATA_WIDTH-1:0] node_194;
    wire [DATA_WIDTH-1:0] node_195;
    wire [DATA_WIDTH-1:0] node_196;
    wire [DATA_WIDTH-1:0] node_197;
    wire [DATA_WIDTH-1:0] node_198;
    wire [DATA_WIDTH-1:0] node_199;
    wire [DATA_WIDTH-1:0] node_200;
    wire [DATA_WIDTH-1:0] node_201;
    wire [DATA_WIDTH-1:0] node_202;
    wire [DATA_WIDTH-1:0] node_203;
    wire [DATA_WIDTH-1:0] node_204;
    wire [DATA_WIDTH-1:0] node_205;
    wire [DATA_WIDTH-1:0] node_206;
    wire [DATA_WIDTH-1:0] node_207;
    wire [DATA_WIDTH-1:0] node_208;
    wire [DATA_WIDTH-1:0] node_209;
    wire [DATA_WIDTH-1:0] node_210;
    wire [DATA_WIDTH-1:0] node_211;
    wire [DATA_WIDTH-1:0] node_212;
    wire [DATA_WIDTH-1:0] node_213;
    wire [DATA_WIDTH-1:0] node_214;
    wire [DATA_WIDTH-1:0] node_215;
    wire [DATA_WIDTH-1:0] node_216;
    wire [DATA_WIDTH-1:0] node_217;
    wire [DATA_WIDTH-1:0] node_218;
    wire [DATA_WIDTH-1:0] node_219;
    wire [DATA_WIDTH-1:0] node_220;
    wire [DATA_WIDTH-1:0] node_221;
    wire [DATA_WIDTH-1:0] node_222;
    wire [DATA_WIDTH-1:0] node_223;
    wire [DATA_WIDTH-1:0] node_224;
    wire [DATA_WIDTH-1:0] node_225;
    wire [DATA_WIDTH-1:0] node_226;
    wire [DATA_WIDTH-1:0] node_227;
    wire [DATA_WIDTH-1:0] node_228;
    wire [DATA_WIDTH-1:0] node_229;
    wire [DATA_WIDTH-1:0] node_230;
    wire [DATA_WIDTH-1:0] node_231;
    wire [DATA_WIDTH-1:0] node_232;
    wire [DATA_WIDTH-1:0] node_233;
    wire [DATA_WIDTH-1:0] node_234;
    wire [DATA_WIDTH-1:0] node_235;
    wire [DATA_WIDTH-1:0] node_236;
    wire [DATA_WIDTH-1:0] node_237;
    wire [DATA_WIDTH-1:0] node_238;
    wire [DATA_WIDTH-1:0] node_239;
    wire [DATA_WIDTH-1:0] node_240;
    wire [DATA_WIDTH-1:0] node_241;
    wire [DATA_WIDTH-1:0] node_242;
    wire [DATA_WIDTH-1:0] node_243;
    wire [DATA_WIDTH-1:0] node_244;
    wire [DATA_WIDTH-1:0] node_245;
    wire [DATA_WIDTH-1:0] node_246;
    wire [DATA_WIDTH-1:0] node_247;
    wire [DATA_WIDTH-1:0] node_248;
    wire [DATA_WIDTH-1:0] node_249;
    wire [DATA_WIDTH-1:0] node_250;
    wire [DATA_WIDTH-1:0] node_251;
    wire [DATA_WIDTH-1:0] node_252;
    wire [DATA_WIDTH-1:0] node_253;
    wire [DATA_WIDTH-1:0] node_254;
    wire [DATA_WIDTH-1:0] node_255;
    wire [DATA_WIDTH-1:0] node_256;
    wire [DATA_WIDTH-1:0] node_257;
    wire [DATA_WIDTH-1:0] node_258;
    wire [DATA_WIDTH-1:0] node_259;
    wire [DATA_WIDTH-1:0] node_260;
    wire [DATA_WIDTH-1:0] node_261;
    wire [DATA_WIDTH-1:0] node_262;
    wire [DATA_WIDTH-1:0] node_263;
    wire [DATA_WIDTH-1:0] node_264;
    wire [DATA_WIDTH-1:0] node_265;
    wire [DATA_WIDTH-1:0] node_266;
    wire [DATA_WIDTH-1:0] node_267;
    wire [DATA_WIDTH-1:0] node_268;
    wire [DATA_WIDTH-1:0] node_269;
    wire [DATA_WIDTH-1:0] node_270;
    wire [DATA_WIDTH-1:0] node_271;
    wire [DATA_WIDTH-1:0] node_272;
    wire [DATA_WIDTH-1:0] node_273;
    wire [DATA_WIDTH-1:0] node_274;
    wire [DATA_WIDTH-1:0] node_275;
    wire [DATA_WIDTH-1:0] node_276;
    wire [DATA_WIDTH-1:0] node_277;
    wire [DATA_WIDTH-1:0] node_278;
    wire [DATA_WIDTH-1:0] node_279;
    wire [DATA_WIDTH-1:0] node_280;
    wire [DATA_WIDTH-1:0] node_281;
    wire [DATA_WIDTH-1:0] node_282;
    wire [DATA_WIDTH-1:0] node_283;
    wire [DATA_WIDTH-1:0] node_284;
    wire [DATA_WIDTH-1:0] node_285;
    wire [DATA_WIDTH-1:0] node_286;
    wire [DATA_WIDTH-1:0] node_287;
    wire [DATA_WIDTH-1:0] node_288;
    wire [DATA_WIDTH-1:0] node_289;
    wire [DATA_WIDTH-1:0] node_290;
    wire [DATA_WIDTH-1:0] node_291;
    wire [DATA_WIDTH-1:0] node_292;
    wire [DATA_WIDTH-1:0] node_293;
    wire [DATA_WIDTH-1:0] node_294;
    wire [DATA_WIDTH-1:0] node_295;
    wire [DATA_WIDTH-1:0] node_296;
    wire [DATA_WIDTH-1:0] node_297;
    wire [DATA_WIDTH-1:0] node_298;
    wire [DATA_WIDTH-1:0] node_299;
    wire [DATA_WIDTH-1:0] node_300;
    wire [DATA_WIDTH-1:0] node_301;
    wire [DATA_WIDTH-1:0] node_302;
    wire [DATA_WIDTH-1:0] node_303;
    wire [DATA_WIDTH-1:0] node_304;
    wire [DATA_WIDTH-1:0] node_305;
    wire [DATA_WIDTH-1:0] node_306;
    wire [DATA_WIDTH-1:0] node_307;
    wire [DATA_WIDTH-1:0] node_308;
    wire [DATA_WIDTH-1:0] node_309;
    wire [DATA_WIDTH-1:0] node_310;
    wire [DATA_WIDTH-1:0] node_311;
    wire [DATA_WIDTH-1:0] node_312;
    wire [DATA_WIDTH-1:0] node_313;
    wire [DATA_WIDTH-1:0] node_314;
    wire [DATA_WIDTH-1:0] node_315;
    wire [DATA_WIDTH-1:0] node_316;
    wire [DATA_WIDTH-1:0] node_317;
    wire [DATA_WIDTH-1:0] node_318;
    wire [DATA_WIDTH-1:0] node_319;
    wire [DATA_WIDTH-1:0] node_320;
    wire [DATA_WIDTH-1:0] node_321;
    wire [DATA_WIDTH-1:0] node_322;
    wire [DATA_WIDTH-1:0] node_323;
    wire [DATA_WIDTH-1:0] node_324;
    wire [DATA_WIDTH-1:0] node_325;
    wire [DATA_WIDTH-1:0] node_326;
    wire [DATA_WIDTH-1:0] node_327;
    wire [DATA_WIDTH-1:0] node_328;
    wire [DATA_WIDTH-1:0] node_329;
    wire [DATA_WIDTH-1:0] node_330;
    wire [DATA_WIDTH-1:0] node_331;
    wire [DATA_WIDTH-1:0] node_332;
    wire [DATA_WIDTH-1:0] node_333;
    wire [DATA_WIDTH-1:0] node_334;
    wire [DATA_WIDTH-1:0] node_335;
    wire [DATA_WIDTH-1:0] node_336;
    wire [DATA_WIDTH-1:0] node_337;
    wire [DATA_WIDTH-1:0] node_338;
    wire [DATA_WIDTH-1:0] node_339;
    wire [DATA_WIDTH-1:0] node_340;
    wire [DATA_WIDTH-1:0] node_341;
    wire [DATA_WIDTH-1:0] node_342;
    wire [DATA_WIDTH-1:0] node_343;
    wire [DATA_WIDTH-1:0] node_344;
    wire [DATA_WIDTH-1:0] node_345;
    wire [DATA_WIDTH-1:0] node_346;
    wire [DATA_WIDTH-1:0] node_347;
    wire [DATA_WIDTH-1:0] node_348;
    wire [DATA_WIDTH-1:0] node_349;
    wire [DATA_WIDTH-1:0] node_350;
    wire [DATA_WIDTH-1:0] node_351;
    wire [DATA_WIDTH-1:0] node_352;
    wire [DATA_WIDTH-1:0] node_353;
    wire [DATA_WIDTH-1:0] node_354;
    wire [DATA_WIDTH-1:0] node_355;
    wire [DATA_WIDTH-1:0] node_356;
    wire [DATA_WIDTH-1:0] node_357;
    wire [DATA_WIDTH-1:0] node_358;
    wire [DATA_WIDTH-1:0] node_359;
    wire [DATA_WIDTH-1:0] node_360;
    wire [DATA_WIDTH-1:0] node_361;
    wire [DATA_WIDTH-1:0] node_362;
    wire [DATA_WIDTH-1:0] node_363;
    wire [DATA_WIDTH-1:0] node_364;
    wire [DATA_WIDTH-1:0] node_365;
    wire [DATA_WIDTH-1:0] node_366;
    wire [DATA_WIDTH-1:0] node_367;
    wire [DATA_WIDTH-1:0] node_368;
    wire [DATA_WIDTH-1:0] node_369;
    wire [DATA_WIDTH-1:0] node_370;
    wire [DATA_WIDTH-1:0] node_371;
    wire [DATA_WIDTH-1:0] node_372;
    wire [DATA_WIDTH-1:0] node_373;
    wire [DATA_WIDTH-1:0] node_374;
    wire [DATA_WIDTH-1:0] node_375;
    wire [DATA_WIDTH-1:0] node_376;
    wire [DATA_WIDTH-1:0] node_377;
    wire [DATA_WIDTH-1:0] node_378;
    wire [DATA_WIDTH-1:0] node_379;
    wire [DATA_WIDTH-1:0] node_380;
    wire [DATA_WIDTH-1:0] node_381;
    wire [DATA_WIDTH-1:0] node_382;
    wire [DATA_WIDTH-1:0] node_383;
    wire [DATA_WIDTH-1:0] node_384;
    wire [DATA_WIDTH-1:0] node_385;
    wire [DATA_WIDTH-1:0] node_386;
    wire [DATA_WIDTH-1:0] node_387;
    wire [DATA_WIDTH-1:0] node_388;
    wire [DATA_WIDTH-1:0] node_389;
    wire [DATA_WIDTH-1:0] node_390;
    wire [DATA_WIDTH-1:0] node_391;
    wire [DATA_WIDTH-1:0] node_392;
    wire [DATA_WIDTH-1:0] node_393;
    wire [DATA_WIDTH-1:0] node_394;
    wire [DATA_WIDTH-1:0] node_395;
    wire [DATA_WIDTH-1:0] node_396;
    wire [DATA_WIDTH-1:0] node_397;
    wire [DATA_WIDTH-1:0] node_398;
    wire [DATA_WIDTH-1:0] node_399;
    wire [DATA_WIDTH-1:0] node_400;
    wire [DATA_WIDTH-1:0] node_401;
    wire [DATA_WIDTH-1:0] node_402;
    wire [DATA_WIDTH-1:0] node_403;
    wire [DATA_WIDTH-1:0] node_404;
    wire [DATA_WIDTH-1:0] node_405;
    wire [DATA_WIDTH-1:0] node_406;
    wire [DATA_WIDTH-1:0] node_407;
    wire [DATA_WIDTH-1:0] node_408;
    wire [DATA_WIDTH-1:0] node_409;
    wire [DATA_WIDTH-1:0] node_410;
    wire [DATA_WIDTH-1:0] node_411;
    wire [DATA_WIDTH-1:0] node_412;
    wire [DATA_WIDTH-1:0] node_413;
    wire [DATA_WIDTH-1:0] node_414;
    wire [DATA_WIDTH-1:0] node_415;
    wire [DATA_WIDTH-1:0] node_416;
    wire [DATA_WIDTH-1:0] node_417;
    wire [DATA_WIDTH-1:0] node_418;
    wire [DATA_WIDTH-1:0] node_419;
    wire [DATA_WIDTH-1:0] node_420;
    wire [DATA_WIDTH-1:0] node_421;
    wire [DATA_WIDTH-1:0] node_422;
    wire [DATA_WIDTH-1:0] node_423;
    wire [DATA_WIDTH-1:0] node_424;
    wire [DATA_WIDTH-1:0] node_425;
    wire [DATA_WIDTH-1:0] node_426;
    wire [DATA_WIDTH-1:0] node_427;
    wire [DATA_WIDTH-1:0] node_428;
    wire [DATA_WIDTH-1:0] node_429;
    wire [DATA_WIDTH-1:0] node_430;
    wire [DATA_WIDTH-1:0] node_431;
    wire [DATA_WIDTH-1:0] node_432;
    wire [DATA_WIDTH-1:0] node_433;
    wire [DATA_WIDTH-1:0] node_434;
    wire [DATA_WIDTH-1:0] node_435;
    wire [DATA_WIDTH-1:0] node_436;
    wire [DATA_WIDTH-1:0] node_437;
    wire [DATA_WIDTH-1:0] node_438;
    wire [DATA_WIDTH-1:0] node_439;
    wire [DATA_WIDTH-1:0] node_440;
    wire [DATA_WIDTH-1:0] node_441;
    wire [DATA_WIDTH-1:0] node_442;
    wire [DATA_WIDTH-1:0] node_443;
    wire [DATA_WIDTH-1:0] node_444;
    wire [DATA_WIDTH-1:0] node_445;
    wire [DATA_WIDTH-1:0] node_446;
    wire [DATA_WIDTH-1:0] node_447;
    wire [DATA_WIDTH-1:0] node_448;
    wire [DATA_WIDTH-1:0] node_449;
    wire [DATA_WIDTH-1:0] node_450;
    wire [DATA_WIDTH-1:0] node_451;
    wire [DATA_WIDTH-1:0] node_452;
    wire [DATA_WIDTH-1:0] node_453;
    wire [DATA_WIDTH-1:0] node_454;
    wire [DATA_WIDTH-1:0] node_455;
    wire [DATA_WIDTH-1:0] node_456;
    wire [DATA_WIDTH-1:0] node_457;
    wire [DATA_WIDTH-1:0] node_458;
    wire [DATA_WIDTH-1:0] node_459;
    wire [DATA_WIDTH-1:0] node_460;
    wire [DATA_WIDTH-1:0] node_461;
    wire [DATA_WIDTH-1:0] node_462;
    wire [DATA_WIDTH-1:0] node_463;
    wire [DATA_WIDTH-1:0] node_464;
    wire [DATA_WIDTH-1:0] node_465;
    wire [DATA_WIDTH-1:0] node_466;
    wire [DATA_WIDTH-1:0] node_467;
    wire [DATA_WIDTH-1:0] node_468;
    wire [DATA_WIDTH-1:0] node_469;
    wire [DATA_WIDTH-1:0] node_470;
    wire [DATA_WIDTH-1:0] node_471;
    wire [DATA_WIDTH-1:0] node_472;
    wire [DATA_WIDTH-1:0] node_473;
    wire [DATA_WIDTH-1:0] node_474;
    wire [DATA_WIDTH-1:0] node_475;
    wire [DATA_WIDTH-1:0] node_476;
    wire [DATA_WIDTH-1:0] node_477;
    wire [DATA_WIDTH-1:0] node_478;
    wire [DATA_WIDTH-1:0] node_479;
    wire [DATA_WIDTH-1:0] node_480;
    wire [DATA_WIDTH-1:0] node_481;
    wire [DATA_WIDTH-1:0] node_482;
    wire [DATA_WIDTH-1:0] node_483;
    wire [DATA_WIDTH-1:0] node_484;
    wire [DATA_WIDTH-1:0] node_485;
    wire [DATA_WIDTH-1:0] node_486;
    wire [DATA_WIDTH-1:0] node_487;
    wire [DATA_WIDTH-1:0] node_488;
    wire [DATA_WIDTH-1:0] node_489;
    wire [DATA_WIDTH-1:0] node_490;
    wire [DATA_WIDTH-1:0] node_491;
    wire [DATA_WIDTH-1:0] node_492;
    wire [DATA_WIDTH-1:0] node_493;
    wire [DATA_WIDTH-1:0] node_494;
    wire [DATA_WIDTH-1:0] node_495;
    wire [DATA_WIDTH-1:0] node_496;
    wire [DATA_WIDTH-1:0] node_497;
    wire [DATA_WIDTH-1:0] node_498;
    wire [DATA_WIDTH-1:0] node_499;
    wire [DATA_WIDTH-1:0] node_500;
    wire [DATA_WIDTH-1:0] node_501;
    wire [DATA_WIDTH-1:0] node_502;
    wire [DATA_WIDTH-1:0] node_503;
    wire [DATA_WIDTH-1:0] node_504;
    wire [DATA_WIDTH-1:0] node_505;
    wire [DATA_WIDTH-1:0] node_506;
    wire [DATA_WIDTH-1:0] node_507;
    wire [DATA_WIDTH-1:0] node_508;
    wire [DATA_WIDTH-1:0] node_509;
    wire [DATA_WIDTH-1:0] node_510;
    wire [DATA_WIDTH-1:0] node_511;
    wire [DATA_WIDTH-1:0] node_512;
    wire [DATA_WIDTH-1:0] node_513;
    wire [DATA_WIDTH-1:0] node_514;
    wire [DATA_WIDTH-1:0] node_515;
    wire [DATA_WIDTH-1:0] node_516;
    wire [DATA_WIDTH-1:0] node_517;
    wire [DATA_WIDTH-1:0] node_518;
    wire [DATA_WIDTH-1:0] node_519;
    wire [DATA_WIDTH-1:0] node_520;
    wire [DATA_WIDTH-1:0] node_521;
    wire [DATA_WIDTH-1:0] node_522;
    wire [DATA_WIDTH-1:0] node_523;
    wire [DATA_WIDTH-1:0] node_524;
    wire [DATA_WIDTH-1:0] node_525;
    wire [DATA_WIDTH-1:0] node_526;
    wire [DATA_WIDTH-1:0] node_527;
    wire [DATA_WIDTH-1:0] node_528;
    wire [DATA_WIDTH-1:0] node_529;
    wire [DATA_WIDTH-1:0] node_530;
    wire [DATA_WIDTH-1:0] node_531;
    wire [DATA_WIDTH-1:0] node_532;
    wire [DATA_WIDTH-1:0] node_533;
    wire [DATA_WIDTH-1:0] node_534;
    wire [DATA_WIDTH-1:0] node_535;
    wire [DATA_WIDTH-1:0] node_536;
    wire [DATA_WIDTH-1:0] node_537;
    wire [DATA_WIDTH-1:0] node_538;
    wire [DATA_WIDTH-1:0] node_539;
    wire [DATA_WIDTH-1:0] node_540;
    wire [DATA_WIDTH-1:0] node_541;
    wire [DATA_WIDTH-1:0] node_542;
    wire [DATA_WIDTH-1:0] node_543;
    wire [DATA_WIDTH-1:0] node_544;
    wire [DATA_WIDTH-1:0] node_545;
    wire [DATA_WIDTH-1:0] node_546;
    wire [DATA_WIDTH-1:0] node_547;
    wire [DATA_WIDTH-1:0] node_548;
    wire [DATA_WIDTH-1:0] node_549;
    wire [DATA_WIDTH-1:0] node_550;
    wire [DATA_WIDTH-1:0] node_551;
    wire [DATA_WIDTH-1:0] node_552;
    wire [DATA_WIDTH-1:0] node_553;
    wire [DATA_WIDTH-1:0] node_554;
    wire [DATA_WIDTH-1:0] node_555;
    wire [DATA_WIDTH-1:0] node_556;
    wire [DATA_WIDTH-1:0] node_557;
    wire [DATA_WIDTH-1:0] node_558;
    wire [DATA_WIDTH-1:0] node_559;
    wire [DATA_WIDTH-1:0] node_560;
    wire [DATA_WIDTH-1:0] node_561;
    wire [DATA_WIDTH-1:0] node_562;
    wire [DATA_WIDTH-1:0] node_563;
    wire [DATA_WIDTH-1:0] node_564;
    wire [DATA_WIDTH-1:0] node_565;
    wire [DATA_WIDTH-1:0] node_566;
    wire [DATA_WIDTH-1:0] node_567;
    wire [DATA_WIDTH-1:0] node_568;
    wire [DATA_WIDTH-1:0] node_569;
    wire [DATA_WIDTH-1:0] node_570;
    wire [DATA_WIDTH-1:0] node_571;
    wire [DATA_WIDTH-1:0] node_572;
    wire [DATA_WIDTH-1:0] node_573;
    wire [DATA_WIDTH-1:0] node_574;
    wire [DATA_WIDTH-1:0] node_575;
    wire [DATA_WIDTH-1:0] node_576;
    wire [DATA_WIDTH-1:0] node_577;
    wire [DATA_WIDTH-1:0] node_578;
    wire [DATA_WIDTH-1:0] node_579;
    wire [DATA_WIDTH-1:0] node_580;
    wire [DATA_WIDTH-1:0] node_581;
    wire [DATA_WIDTH-1:0] node_582;
    wire [DATA_WIDTH-1:0] node_583;
    wire [DATA_WIDTH-1:0] node_584;
    wire [DATA_WIDTH-1:0] node_585;
    wire [DATA_WIDTH-1:0] node_586;
    wire [DATA_WIDTH-1:0] node_587;
    wire [DATA_WIDTH-1:0] node_588;
    wire [DATA_WIDTH-1:0] node_589;
    wire [DATA_WIDTH-1:0] node_590;
    wire [DATA_WIDTH-1:0] node_591;
    wire [DATA_WIDTH-1:0] node_592;
    wire [DATA_WIDTH-1:0] node_593;
    wire [DATA_WIDTH-1:0] node_594;
    wire [DATA_WIDTH-1:0] node_595;
    wire [DATA_WIDTH-1:0] node_596;
    wire [DATA_WIDTH-1:0] node_597;
    wire [DATA_WIDTH-1:0] node_598;
    wire [DATA_WIDTH-1:0] node_599;
    wire [DATA_WIDTH-1:0] node_600;
    wire [DATA_WIDTH-1:0] node_601;
    wire [DATA_WIDTH-1:0] node_602;
    wire [DATA_WIDTH-1:0] node_603;
    wire [DATA_WIDTH-1:0] node_604;
    wire [DATA_WIDTH-1:0] node_605;
    wire [DATA_WIDTH-1:0] node_606;
    wire [DATA_WIDTH-1:0] node_607;
    wire [DATA_WIDTH-1:0] node_608;
    wire [DATA_WIDTH-1:0] node_609;
    wire [DATA_WIDTH-1:0] node_610;
    wire [DATA_WIDTH-1:0] node_611;
    wire [DATA_WIDTH-1:0] node_612;
    wire [DATA_WIDTH-1:0] node_613;
    wire [DATA_WIDTH-1:0] node_614;
    wire [DATA_WIDTH-1:0] node_615;
    wire [DATA_WIDTH-1:0] node_616;
    wire [DATA_WIDTH-1:0] node_617;
    wire [DATA_WIDTH-1:0] node_618;
    wire [DATA_WIDTH-1:0] node_619;
    wire [DATA_WIDTH-1:0] node_620;
    wire [DATA_WIDTH-1:0] node_621;
    wire [DATA_WIDTH-1:0] node_622;
    wire [DATA_WIDTH-1:0] node_623;
    wire [DATA_WIDTH-1:0] node_624;
    wire [DATA_WIDTH-1:0] node_625;
    wire [DATA_WIDTH-1:0] node_626;
    wire [DATA_WIDTH-1:0] node_627;
    wire [DATA_WIDTH-1:0] node_628;
    wire [DATA_WIDTH-1:0] node_629;
    wire [DATA_WIDTH-1:0] node_630;
    wire [DATA_WIDTH-1:0] node_631;
    wire [DATA_WIDTH-1:0] node_632;
    wire [DATA_WIDTH-1:0] node_633;
    wire [DATA_WIDTH-1:0] node_634;
    wire [DATA_WIDTH-1:0] node_635;
    wire [DATA_WIDTH-1:0] node_636;
    wire [DATA_WIDTH-1:0] node_637;
    wire [DATA_WIDTH-1:0] node_638;
    wire [DATA_WIDTH-1:0] node_639;
    wire [DATA_WIDTH-1:0] node_640;
    wire [DATA_WIDTH-1:0] node_641;
    wire [DATA_WIDTH-1:0] node_642;
    wire [DATA_WIDTH-1:0] node_643;
    wire [DATA_WIDTH-1:0] node_644;
    wire [DATA_WIDTH-1:0] node_645;
    wire [DATA_WIDTH-1:0] node_646;
    wire [DATA_WIDTH-1:0] node_647;
    wire [DATA_WIDTH-1:0] node_648;
    wire [DATA_WIDTH-1:0] node_649;
    wire [DATA_WIDTH-1:0] node_650;
    wire [DATA_WIDTH-1:0] node_651;
    wire [DATA_WIDTH-1:0] node_652;
    wire [DATA_WIDTH-1:0] node_653;
    wire [DATA_WIDTH-1:0] node_654;
    wire [DATA_WIDTH-1:0] node_655;
    wire [DATA_WIDTH-1:0] node_656;
    wire [DATA_WIDTH-1:0] node_657;
    wire [DATA_WIDTH-1:0] node_658;
    wire [DATA_WIDTH-1:0] node_659;
    wire [DATA_WIDTH-1:0] node_660;
    wire [DATA_WIDTH-1:0] node_661;
    wire [DATA_WIDTH-1:0] node_662;
    wire [DATA_WIDTH-1:0] node_663;
    wire [DATA_WIDTH-1:0] node_664;
    wire [DATA_WIDTH-1:0] node_665;
    wire [DATA_WIDTH-1:0] node_666;
    wire [DATA_WIDTH-1:0] node_667;
    wire [DATA_WIDTH-1:0] node_668;
    wire [DATA_WIDTH-1:0] node_669;
    wire [DATA_WIDTH-1:0] node_670;
    wire [DATA_WIDTH-1:0] node_671;
    wire [DATA_WIDTH-1:0] node_672;
    wire [DATA_WIDTH-1:0] node_673;
    wire [DATA_WIDTH-1:0] node_674;
    wire [DATA_WIDTH-1:0] node_675;
    wire [DATA_WIDTH-1:0] node_676;
    wire [DATA_WIDTH-1:0] node_677;
    wire [DATA_WIDTH-1:0] node_678;
    wire [DATA_WIDTH-1:0] node_679;
    wire [DATA_WIDTH-1:0] node_680;
    wire [DATA_WIDTH-1:0] node_681;
    wire [DATA_WIDTH-1:0] node_682;
    wire [DATA_WIDTH-1:0] node_683;
    wire [DATA_WIDTH-1:0] node_684;
    wire [DATA_WIDTH-1:0] node_685;
    wire [DATA_WIDTH-1:0] node_686;
    wire [DATA_WIDTH-1:0] node_687;
    wire [DATA_WIDTH-1:0] node_688;
    wire [DATA_WIDTH-1:0] node_689;
    wire [DATA_WIDTH-1:0] node_690;
    wire [DATA_WIDTH-1:0] node_691;
    wire [DATA_WIDTH-1:0] node_692;
    wire [DATA_WIDTH-1:0] node_693;
    wire [DATA_WIDTH-1:0] node_694;
    wire [DATA_WIDTH-1:0] node_695;
    wire [DATA_WIDTH-1:0] node_696;
    wire [DATA_WIDTH-1:0] node_697;
    wire [DATA_WIDTH-1:0] node_698;
    wire [DATA_WIDTH-1:0] node_699;
    wire [DATA_WIDTH-1:0] node_700;
    wire [DATA_WIDTH-1:0] node_701;
    wire [DATA_WIDTH-1:0] node_702;
    wire [DATA_WIDTH-1:0] node_703;
    wire [DATA_WIDTH-1:0] node_704;
    wire [DATA_WIDTH-1:0] node_705;
    wire [DATA_WIDTH-1:0] node_706;
    wire [DATA_WIDTH-1:0] node_707;
    wire [DATA_WIDTH-1:0] node_708;
    wire [DATA_WIDTH-1:0] node_709;
    wire [DATA_WIDTH-1:0] node_710;
    wire [DATA_WIDTH-1:0] node_711;
    wire [DATA_WIDTH-1:0] node_712;
    wire [DATA_WIDTH-1:0] node_713;
    wire [DATA_WIDTH-1:0] node_714;
    wire [DATA_WIDTH-1:0] node_715;
    wire [DATA_WIDTH-1:0] node_716;
    wire [DATA_WIDTH-1:0] node_717;
    wire [DATA_WIDTH-1:0] node_718;
    wire [DATA_WIDTH-1:0] node_719;
    wire [DATA_WIDTH-1:0] node_720;
    wire [DATA_WIDTH-1:0] node_721;
    wire [DATA_WIDTH-1:0] node_722;
    wire [DATA_WIDTH-1:0] node_723;
    wire [DATA_WIDTH-1:0] node_724;
    wire [DATA_WIDTH-1:0] node_725;
    wire [DATA_WIDTH-1:0] node_726;
    wire [DATA_WIDTH-1:0] node_727;
    wire [DATA_WIDTH-1:0] node_728;
    wire [DATA_WIDTH-1:0] node_729;
    wire [DATA_WIDTH-1:0] node_730;
    wire [DATA_WIDTH-1:0] node_731;
    wire [DATA_WIDTH-1:0] node_732;
    wire [DATA_WIDTH-1:0] node_733;
    wire [DATA_WIDTH-1:0] node_734;
    wire [DATA_WIDTH-1:0] node_735;
    wire [DATA_WIDTH-1:0] node_736;
    wire [DATA_WIDTH-1:0] node_737;
    wire [DATA_WIDTH-1:0] node_738;
    wire [DATA_WIDTH-1:0] node_739;
    wire [DATA_WIDTH-1:0] node_740;
    wire [DATA_WIDTH-1:0] node_741;
    wire [DATA_WIDTH-1:0] node_742;
    wire [DATA_WIDTH-1:0] node_743;
    wire [DATA_WIDTH-1:0] node_744;
    wire [DATA_WIDTH-1:0] node_745;
    wire [DATA_WIDTH-1:0] node_746;
    wire [DATA_WIDTH-1:0] node_747;
    wire [DATA_WIDTH-1:0] node_748;
    wire [DATA_WIDTH-1:0] node_749;
    wire [DATA_WIDTH-1:0] node_750;
    wire [DATA_WIDTH-1:0] node_751;
    wire [DATA_WIDTH-1:0] node_752;
    wire [DATA_WIDTH-1:0] node_753;
    wire [DATA_WIDTH-1:0] node_754;
    wire [DATA_WIDTH-1:0] node_755;
    wire [DATA_WIDTH-1:0] node_756;
    wire [DATA_WIDTH-1:0] node_757;
    wire [DATA_WIDTH-1:0] node_758;
    wire [DATA_WIDTH-1:0] node_759;
    wire [DATA_WIDTH-1:0] node_760;
    wire [DATA_WIDTH-1:0] node_761;
    wire [DATA_WIDTH-1:0] node_762;
    wire [DATA_WIDTH-1:0] node_763;
    wire [DATA_WIDTH-1:0] node_764;
    wire [DATA_WIDTH-1:0] node_765;
    wire [DATA_WIDTH-1:0] node_766;
    wire [DATA_WIDTH-1:0] node_767;
    wire [DATA_WIDTH-1:0] node_768;
    wire [DATA_WIDTH-1:0] node_769;
    wire [DATA_WIDTH-1:0] node_770;
    wire [DATA_WIDTH-1:0] node_771;
    wire [DATA_WIDTH-1:0] node_772;
    wire [DATA_WIDTH-1:0] node_773;
    wire [DATA_WIDTH-1:0] node_774;
    wire [DATA_WIDTH-1:0] node_775;
    wire [DATA_WIDTH-1:0] node_776;
    wire [DATA_WIDTH-1:0] node_777;
    wire [DATA_WIDTH-1:0] node_778;
    wire [DATA_WIDTH-1:0] node_779;
    wire [DATA_WIDTH-1:0] node_780;
    wire [DATA_WIDTH-1:0] node_781;
    wire [DATA_WIDTH-1:0] node_782;
    wire [DATA_WIDTH-1:0] node_783;
    wire [DATA_WIDTH-1:0] node_784;
    wire [DATA_WIDTH-1:0] node_785;
    wire [DATA_WIDTH-1:0] node_786;
    wire [DATA_WIDTH-1:0] node_787;
    wire [DATA_WIDTH-1:0] node_788;
    wire [DATA_WIDTH-1:0] node_789;
    wire [DATA_WIDTH-1:0] node_790;
    wire [DATA_WIDTH-1:0] node_791;
    wire [DATA_WIDTH-1:0] node_792;
    wire [DATA_WIDTH-1:0] node_793;
    wire [DATA_WIDTH-1:0] node_794;
    wire [DATA_WIDTH-1:0] node_795;
    wire [DATA_WIDTH-1:0] node_796;
    wire [DATA_WIDTH-1:0] node_797;
    wire [DATA_WIDTH-1:0] node_798;
    wire [DATA_WIDTH-1:0] node_799;
    wire [DATA_WIDTH-1:0] node_800;
    wire [DATA_WIDTH-1:0] node_801;
    wire [DATA_WIDTH-1:0] node_802;
    wire [DATA_WIDTH-1:0] node_803;
    wire [DATA_WIDTH-1:0] node_804;
    wire [DATA_WIDTH-1:0] node_805;
    wire [DATA_WIDTH-1:0] node_806;
    wire [DATA_WIDTH-1:0] node_807;
    wire [DATA_WIDTH-1:0] node_808;
    wire [DATA_WIDTH-1:0] node_809;
    wire [DATA_WIDTH-1:0] node_810;
    wire [DATA_WIDTH-1:0] node_811;
    wire [DATA_WIDTH-1:0] node_812;
    wire [DATA_WIDTH-1:0] node_813;
    wire [DATA_WIDTH-1:0] node_814;
    wire [DATA_WIDTH-1:0] node_815;
    wire [DATA_WIDTH-1:0] node_816;
    wire [DATA_WIDTH-1:0] node_817;
    wire [DATA_WIDTH-1:0] node_818;
    wire [DATA_WIDTH-1:0] node_819;
    wire [DATA_WIDTH-1:0] node_820;
    wire [DATA_WIDTH-1:0] node_821;
    wire [DATA_WIDTH-1:0] node_822;
    wire [DATA_WIDTH-1:0] node_823;
    wire [DATA_WIDTH-1:0] node_824;
    wire [DATA_WIDTH-1:0] node_825;
    wire [DATA_WIDTH-1:0] node_826;
    wire [DATA_WIDTH-1:0] node_827;
    wire [DATA_WIDTH-1:0] node_828;
    wire [DATA_WIDTH-1:0] node_829;
    wire [DATA_WIDTH-1:0] node_830;
    wire [DATA_WIDTH-1:0] node_831;
    wire [DATA_WIDTH-1:0] node_832;
    wire [DATA_WIDTH-1:0] node_833;
    wire [DATA_WIDTH-1:0] node_834;
    wire [DATA_WIDTH-1:0] node_835;
    wire [DATA_WIDTH-1:0] node_836;
    wire [DATA_WIDTH-1:0] node_837;
    wire [DATA_WIDTH-1:0] node_838;
    wire [DATA_WIDTH-1:0] node_839;
    wire [DATA_WIDTH-1:0] node_840;
    wire [DATA_WIDTH-1:0] node_841;
    wire [DATA_WIDTH-1:0] node_842;
    wire [DATA_WIDTH-1:0] node_843;
    wire [DATA_WIDTH-1:0] node_844;
    wire [DATA_WIDTH-1:0] node_845;
    wire [DATA_WIDTH-1:0] node_846;
    wire [DATA_WIDTH-1:0] node_847;
    wire [DATA_WIDTH-1:0] node_848;
    wire [DATA_WIDTH-1:0] node_849;
    wire [DATA_WIDTH-1:0] node_850;
    wire [DATA_WIDTH-1:0] node_851;
    wire [DATA_WIDTH-1:0] node_852;
    wire [DATA_WIDTH-1:0] node_853;
    wire [DATA_WIDTH-1:0] node_854;
    wire [DATA_WIDTH-1:0] node_855;
    wire [DATA_WIDTH-1:0] node_856;
    wire [DATA_WIDTH-1:0] node_857;
    wire [DATA_WIDTH-1:0] node_858;
    wire [DATA_WIDTH-1:0] node_859;
    wire [DATA_WIDTH-1:0] node_860;
    wire [DATA_WIDTH-1:0] node_861;
    wire [DATA_WIDTH-1:0] node_862;
    wire [DATA_WIDTH-1:0] node_863;
    wire [DATA_WIDTH-1:0] node_864;
    wire [DATA_WIDTH-1:0] node_865;
    wire [DATA_WIDTH-1:0] node_866;
    wire [DATA_WIDTH-1:0] node_867;
    wire [DATA_WIDTH-1:0] node_868;
    wire [DATA_WIDTH-1:0] node_869;
    wire [DATA_WIDTH-1:0] node_870;
    wire [DATA_WIDTH-1:0] node_871;
    wire [DATA_WIDTH-1:0] node_872;
    wire [DATA_WIDTH-1:0] node_873;
    wire [DATA_WIDTH-1:0] node_874;
    wire [DATA_WIDTH-1:0] node_875;
    wire [DATA_WIDTH-1:0] node_876;
    wire [DATA_WIDTH-1:0] node_877;
    wire [DATA_WIDTH-1:0] node_878;
    wire [DATA_WIDTH-1:0] node_879;
    wire [DATA_WIDTH-1:0] node_880;
    wire [DATA_WIDTH-1:0] node_881;
    wire [DATA_WIDTH-1:0] node_882;
    wire [DATA_WIDTH-1:0] node_883;
    wire [DATA_WIDTH-1:0] node_884;
    wire [DATA_WIDTH-1:0] node_885;
    wire [DATA_WIDTH-1:0] node_886;
    wire [DATA_WIDTH-1:0] node_887;
    wire [DATA_WIDTH-1:0] node_888;
    wire [DATA_WIDTH-1:0] node_889;
    wire [DATA_WIDTH-1:0] node_890;
    wire [DATA_WIDTH-1:0] node_891;
    wire [DATA_WIDTH-1:0] node_892;
    wire [DATA_WIDTH-1:0] node_893;
    wire [DATA_WIDTH-1:0] node_894;
    wire [DATA_WIDTH-1:0] node_895;
    wire [DATA_WIDTH-1:0] node_896;
    wire [DATA_WIDTH-1:0] node_897;
    wire [DATA_WIDTH-1:0] node_898;
    wire [DATA_WIDTH-1:0] node_899;
    wire [DATA_WIDTH-1:0] node_900;
    wire [DATA_WIDTH-1:0] node_901;
    wire [DATA_WIDTH-1:0] node_902;
    wire [DATA_WIDTH-1:0] node_903;
    wire [DATA_WIDTH-1:0] node_904;
    wire [DATA_WIDTH-1:0] node_905;
    wire [DATA_WIDTH-1:0] node_906;
    wire [DATA_WIDTH-1:0] node_907;
    wire [DATA_WIDTH-1:0] node_908;
    wire [DATA_WIDTH-1:0] node_909;
    wire [DATA_WIDTH-1:0] node_910;
    wire [DATA_WIDTH-1:0] node_911;
    wire [DATA_WIDTH-1:0] node_912;
    wire [DATA_WIDTH-1:0] node_913;
    wire [DATA_WIDTH-1:0] node_914;
    wire [DATA_WIDTH-1:0] node_915;
    wire [DATA_WIDTH-1:0] node_916;
    wire [DATA_WIDTH-1:0] node_917;
    wire [DATA_WIDTH-1:0] node_918;
    wire [DATA_WIDTH-1:0] node_919;
    wire [DATA_WIDTH-1:0] node_920;
    wire [DATA_WIDTH-1:0] node_921;
    wire [DATA_WIDTH-1:0] node_922;
    wire [DATA_WIDTH-1:0] node_923;
    wire [DATA_WIDTH-1:0] node_924;
    wire [DATA_WIDTH-1:0] node_925;
    wire [DATA_WIDTH-1:0] node_926;
    wire [DATA_WIDTH-1:0] node_927;
    wire [DATA_WIDTH-1:0] node_928;
    wire [DATA_WIDTH-1:0] node_929;
    wire [DATA_WIDTH-1:0] node_930;
    wire [DATA_WIDTH-1:0] node_931;
    wire [DATA_WIDTH-1:0] node_932;
    wire [DATA_WIDTH-1:0] node_933;
    wire [DATA_WIDTH-1:0] node_934;
    wire [DATA_WIDTH-1:0] node_935;
    wire [DATA_WIDTH-1:0] node_936;
    wire [DATA_WIDTH-1:0] node_937;
    wire [DATA_WIDTH-1:0] node_938;
    wire [DATA_WIDTH-1:0] node_939;
    wire [DATA_WIDTH-1:0] node_940;
    wire [DATA_WIDTH-1:0] node_941;
    wire [DATA_WIDTH-1:0] node_942;
    wire [DATA_WIDTH-1:0] node_943;
    wire [DATA_WIDTH-1:0] node_944;
    wire [DATA_WIDTH-1:0] node_945;
    wire [DATA_WIDTH-1:0] node_946;
    wire [DATA_WIDTH-1:0] node_947;
    wire [DATA_WIDTH-1:0] node_948;
    wire [DATA_WIDTH-1:0] node_949;
    wire [DATA_WIDTH-1:0] node_950;
    wire [DATA_WIDTH-1:0] node_951;
    wire [DATA_WIDTH-1:0] node_952;
    wire [DATA_WIDTH-1:0] node_953;
    wire [DATA_WIDTH-1:0] node_954;
    wire [DATA_WIDTH-1:0] node_955;
    wire [DATA_WIDTH-1:0] node_956;
    wire [DATA_WIDTH-1:0] node_957;
    wire [DATA_WIDTH-1:0] node_958;
    wire [DATA_WIDTH-1:0] node_959;
    wire [DATA_WIDTH-1:0] node_960;
    wire [DATA_WIDTH-1:0] node_961;
    wire [DATA_WIDTH-1:0] node_962;
    wire [DATA_WIDTH-1:0] node_963;
    wire [DATA_WIDTH-1:0] node_964;
    wire [DATA_WIDTH-1:0] node_965;
    wire [DATA_WIDTH-1:0] node_966;
    wire [DATA_WIDTH-1:0] node_967;
    wire [DATA_WIDTH-1:0] node_968;
    wire [DATA_WIDTH-1:0] node_969;
    wire [DATA_WIDTH-1:0] node_970;
    wire [DATA_WIDTH-1:0] node_971;
    wire [DATA_WIDTH-1:0] node_972;
    wire [DATA_WIDTH-1:0] node_973;
    wire [DATA_WIDTH-1:0] node_974;
    wire [DATA_WIDTH-1:0] node_975;
    wire [DATA_WIDTH-1:0] node_976;
    wire [DATA_WIDTH-1:0] node_977;
    wire [DATA_WIDTH-1:0] node_978;
    wire [DATA_WIDTH-1:0] node_979;
    wire [DATA_WIDTH-1:0] node_980;
    wire [DATA_WIDTH-1:0] node_981;
    wire [DATA_WIDTH-1:0] node_982;
    wire [DATA_WIDTH-1:0] node_983;
    wire [DATA_WIDTH-1:0] node_984;
    wire [DATA_WIDTH-1:0] node_985;
    wire [DATA_WIDTH-1:0] node_986;
    wire [DATA_WIDTH-1:0] node_987;
    wire [DATA_WIDTH-1:0] node_988;
    wire [DATA_WIDTH-1:0] node_989;
    wire [DATA_WIDTH-1:0] node_990;
    wire [DATA_WIDTH-1:0] node_991;
    wire [DATA_WIDTH-1:0] node_992;
    wire [DATA_WIDTH-1:0] node_993;
    wire [DATA_WIDTH-1:0] node_994;
    wire [DATA_WIDTH-1:0] node_995;
    wire [DATA_WIDTH-1:0] node_996;
    wire [DATA_WIDTH-1:0] node_997;
    wire [DATA_WIDTH-1:0] node_998;
    wire [DATA_WIDTH-1:0] node_999;
    wire [DATA_WIDTH-1:0] node_1000;
    wire [DATA_WIDTH-1:0] node_1001;
    wire [DATA_WIDTH-1:0] node_1002;
    wire [DATA_WIDTH-1:0] node_1003;
    wire [DATA_WIDTH-1:0] node_1004;
    wire [DATA_WIDTH-1:0] node_1005;
    wire [DATA_WIDTH-1:0] node_1006;
    wire [DATA_WIDTH-1:0] node_1007;
    wire [DATA_WIDTH-1:0] node_1008;
    wire [DATA_WIDTH-1:0] node_1009;
    wire [DATA_WIDTH-1:0] node_1010;
    wire [DATA_WIDTH-1:0] node_1011;
    wire [DATA_WIDTH-1:0] node_1012;
    wire [DATA_WIDTH-1:0] node_1013;
    wire [DATA_WIDTH-1:0] node_1014;
    wire [DATA_WIDTH-1:0] node_1015;
    wire [DATA_WIDTH-1:0] node_1016;
    wire [DATA_WIDTH-1:0] node_1017;
    wire [DATA_WIDTH-1:0] node_1018;
    wire [DATA_WIDTH-1:0] node_1019;
    wire [DATA_WIDTH-1:0] node_1020;
    wire [DATA_WIDTH-1:0] node_1021;
    wire [DATA_WIDTH-1:0] node_1022;
    wire [DATA_WIDTH-1:0] node_1023;
    wire [DATA_WIDTH-1:0] node_1024;
    wire [DATA_WIDTH-1:0] node_1025;
    wire [DATA_WIDTH-1:0] node_1026;
    wire [DATA_WIDTH-1:0] node_1027;
    wire [DATA_WIDTH-1:0] node_1028;
    wire [DATA_WIDTH-1:0] node_1029;
    wire [DATA_WIDTH-1:0] node_1030;
    wire [DATA_WIDTH-1:0] node_1031;
    wire [DATA_WIDTH-1:0] node_1032;
    wire [DATA_WIDTH-1:0] node_1033;
    wire [DATA_WIDTH-1:0] node_1034;
    wire [DATA_WIDTH-1:0] node_1035;
    wire [DATA_WIDTH-1:0] node_1036;
    wire [DATA_WIDTH-1:0] node_1037;
    wire [DATA_WIDTH-1:0] node_1038;
    wire [DATA_WIDTH-1:0] node_1039;
    wire [DATA_WIDTH-1:0] node_1040;
    wire [DATA_WIDTH-1:0] node_1041;
    wire [DATA_WIDTH-1:0] node_1042;
    wire [DATA_WIDTH-1:0] node_1043;
    wire [DATA_WIDTH-1:0] node_1044;
    wire [DATA_WIDTH-1:0] node_1045;
    wire [DATA_WIDTH-1:0] node_1046;
    wire [DATA_WIDTH-1:0] node_1047;
    wire [DATA_WIDTH-1:0] node_1048;
    wire [DATA_WIDTH-1:0] node_1049;
    wire [DATA_WIDTH-1:0] node_1050;
    wire [DATA_WIDTH-1:0] node_1051;
    wire [DATA_WIDTH-1:0] node_1052;
    wire [DATA_WIDTH-1:0] node_1053;
    wire [DATA_WIDTH-1:0] node_1054;
    wire [DATA_WIDTH-1:0] node_1055;
    wire [DATA_WIDTH-1:0] node_1056;
    wire [DATA_WIDTH-1:0] node_1057;
    wire [DATA_WIDTH-1:0] node_1058;
    wire [DATA_WIDTH-1:0] node_1059;
    wire [DATA_WIDTH-1:0] node_1060;
    wire [DATA_WIDTH-1:0] node_1061;
    wire [DATA_WIDTH-1:0] node_1062;
    wire [DATA_WIDTH-1:0] node_1063;
    wire [DATA_WIDTH-1:0] node_1064;
    wire [DATA_WIDTH-1:0] node_1065;
    wire [DATA_WIDTH-1:0] node_1066;
    wire [DATA_WIDTH-1:0] node_1067;
    wire [DATA_WIDTH-1:0] node_1068;
    wire [DATA_WIDTH-1:0] node_1069;
    wire [DATA_WIDTH-1:0] node_1070;
    wire [DATA_WIDTH-1:0] node_1071;
    wire [DATA_WIDTH-1:0] node_1072;
    wire [DATA_WIDTH-1:0] node_1073;
    wire [DATA_WIDTH-1:0] node_1074;
    wire [DATA_WIDTH-1:0] node_1075;
    wire [DATA_WIDTH-1:0] node_1076;
    wire [DATA_WIDTH-1:0] node_1077;
    wire [DATA_WIDTH-1:0] node_1078;
    wire [DATA_WIDTH-1:0] node_1079;
    wire [DATA_WIDTH-1:0] node_1080;
    wire [DATA_WIDTH-1:0] node_1081;
    wire [DATA_WIDTH-1:0] node_1082;
    wire [DATA_WIDTH-1:0] node_1083;
    wire [DATA_WIDTH-1:0] node_1084;
    wire [DATA_WIDTH-1:0] node_1085;
    wire [DATA_WIDTH-1:0] node_1086;
    wire [DATA_WIDTH-1:0] node_1087;
    wire [DATA_WIDTH-1:0] node_1088;
    wire [DATA_WIDTH-1:0] node_1089;
    wire [DATA_WIDTH-1:0] node_1090;
    wire [DATA_WIDTH-1:0] node_1091;
    wire [DATA_WIDTH-1:0] node_1092;
    wire [DATA_WIDTH-1:0] node_1093;
    wire [DATA_WIDTH-1:0] node_1094;
    wire [DATA_WIDTH-1:0] node_1095;
    wire [DATA_WIDTH-1:0] node_1096;
    wire [DATA_WIDTH-1:0] node_1097;
    wire [DATA_WIDTH-1:0] node_1098;
    wire [DATA_WIDTH-1:0] node_1099;
    wire [DATA_WIDTH-1:0] node_1100;
    wire [DATA_WIDTH-1:0] node_1101;
    wire [DATA_WIDTH-1:0] node_1102;
    wire [DATA_WIDTH-1:0] node_1103;
    wire [DATA_WIDTH-1:0] node_1104;
    wire [DATA_WIDTH-1:0] node_1105;
    wire [DATA_WIDTH-1:0] node_1106;
    wire [DATA_WIDTH-1:0] node_1107;
    wire [DATA_WIDTH-1:0] node_1108;
    wire [DATA_WIDTH-1:0] node_1109;
    wire [DATA_WIDTH-1:0] node_1110;
    wire [DATA_WIDTH-1:0] node_1111;
    wire [DATA_WIDTH-1:0] node_1112;
    wire [DATA_WIDTH-1:0] node_1113;
    wire [DATA_WIDTH-1:0] node_1114;
    wire [DATA_WIDTH-1:0] node_1115;
    wire [DATA_WIDTH-1:0] node_1116;
    wire [DATA_WIDTH-1:0] node_1117;
    wire [DATA_WIDTH-1:0] node_1118;
    wire [DATA_WIDTH-1:0] node_1119;
    wire [DATA_WIDTH-1:0] node_1120;
    wire [DATA_WIDTH-1:0] node_1121;
    wire [DATA_WIDTH-1:0] node_1122;
    wire [DATA_WIDTH-1:0] node_1123;
    wire [DATA_WIDTH-1:0] node_1124;
    wire [DATA_WIDTH-1:0] node_1125;
    wire [DATA_WIDTH-1:0] node_1126;
    wire [DATA_WIDTH-1:0] node_1127;
    wire [DATA_WIDTH-1:0] node_1128;
    wire [DATA_WIDTH-1:0] node_1129;
    wire [DATA_WIDTH-1:0] node_1130;
    wire [DATA_WIDTH-1:0] node_1131;
    wire [DATA_WIDTH-1:0] node_1132;
    wire [DATA_WIDTH-1:0] node_1133;
    wire [DATA_WIDTH-1:0] node_1134;
    wire [DATA_WIDTH-1:0] node_1135;
    wire [DATA_WIDTH-1:0] node_1136;
    wire [DATA_WIDTH-1:0] node_1137;
    wire [DATA_WIDTH-1:0] node_1138;
    wire [DATA_WIDTH-1:0] node_1139;
    wire [DATA_WIDTH-1:0] node_1140;
    wire [DATA_WIDTH-1:0] node_1141;
    wire [DATA_WIDTH-1:0] node_1142;
    wire [DATA_WIDTH-1:0] node_1143;
    wire [DATA_WIDTH-1:0] node_1144;
    wire [DATA_WIDTH-1:0] node_1145;
    wire [DATA_WIDTH-1:0] node_1146;
    wire [DATA_WIDTH-1:0] node_1147;
    wire [DATA_WIDTH-1:0] node_1148;
    wire [DATA_WIDTH-1:0] node_1149;
    wire [DATA_WIDTH-1:0] node_1150;
    wire [DATA_WIDTH-1:0] node_1151;
    wire [DATA_WIDTH-1:0] node_1152;
    wire [DATA_WIDTH-1:0] node_1153;
    wire [DATA_WIDTH-1:0] node_1154;
    wire [DATA_WIDTH-1:0] node_1155;
    wire [DATA_WIDTH-1:0] node_1156;
    wire [DATA_WIDTH-1:0] node_1157;
    wire [DATA_WIDTH-1:0] node_1158;
    wire [DATA_WIDTH-1:0] node_1159;
    wire [DATA_WIDTH-1:0] node_1160;
    wire [DATA_WIDTH-1:0] node_1161;
    wire [DATA_WIDTH-1:0] node_1162;
    wire [DATA_WIDTH-1:0] node_1163;
    wire [DATA_WIDTH-1:0] node_1164;
    wire [DATA_WIDTH-1:0] node_1165;
    wire [DATA_WIDTH-1:0] node_1166;
    wire [DATA_WIDTH-1:0] node_1167;
    wire [DATA_WIDTH-1:0] node_1168;
    wire [DATA_WIDTH-1:0] node_1169;
    wire [DATA_WIDTH-1:0] node_1170;
    wire [DATA_WIDTH-1:0] node_1171;
    wire [DATA_WIDTH-1:0] node_1172;
    wire [DATA_WIDTH-1:0] node_1173;
    wire [DATA_WIDTH-1:0] node_1174;
    wire [DATA_WIDTH-1:0] node_1175;
    wire [DATA_WIDTH-1:0] node_1176;
    wire [DATA_WIDTH-1:0] node_1177;
    wire [DATA_WIDTH-1:0] node_1178;
    wire [DATA_WIDTH-1:0] node_1179;
    wire [DATA_WIDTH-1:0] node_1180;
    wire [DATA_WIDTH-1:0] node_1181;
    wire [DATA_WIDTH-1:0] node_1182;
    wire [DATA_WIDTH-1:0] node_1183;
    wire [DATA_WIDTH-1:0] node_1184;
    wire [DATA_WIDTH-1:0] node_1185;
    wire [DATA_WIDTH-1:0] node_1186;
    wire [DATA_WIDTH-1:0] node_1187;
    wire [DATA_WIDTH-1:0] node_1188;
    wire [DATA_WIDTH-1:0] node_1189;
    wire [DATA_WIDTH-1:0] node_1190;
    wire [DATA_WIDTH-1:0] node_1191;
    wire [DATA_WIDTH-1:0] node_1192;
    wire [DATA_WIDTH-1:0] node_1193;
    wire [DATA_WIDTH-1:0] node_1194;
    wire [DATA_WIDTH-1:0] node_1195;
    wire [DATA_WIDTH-1:0] node_1196;
    wire [DATA_WIDTH-1:0] node_1197;
    wire [DATA_WIDTH-1:0] node_1198;
    wire [DATA_WIDTH-1:0] node_1199;
    wire [DATA_WIDTH-1:0] node_1200;
    wire [DATA_WIDTH-1:0] node_1201;
    wire [DATA_WIDTH-1:0] node_1202;
    wire [DATA_WIDTH-1:0] node_1203;
    wire [DATA_WIDTH-1:0] node_1204;
    wire [DATA_WIDTH-1:0] node_1205;
    wire [DATA_WIDTH-1:0] node_1206;
    wire [DATA_WIDTH-1:0] node_1207;
    wire [DATA_WIDTH-1:0] node_1208;
    wire [DATA_WIDTH-1:0] node_1209;
    wire [DATA_WIDTH-1:0] node_1210;
    wire [DATA_WIDTH-1:0] node_1211;
    wire [DATA_WIDTH-1:0] node_1212;
    wire [DATA_WIDTH-1:0] node_1213;
    wire [DATA_WIDTH-1:0] node_1214;
    wire [DATA_WIDTH-1:0] node_1215;
    wire [DATA_WIDTH-1:0] node_1216;
    wire [DATA_WIDTH-1:0] node_1217;
    wire [DATA_WIDTH-1:0] node_1218;
    wire [DATA_WIDTH-1:0] node_1219;
    wire [DATA_WIDTH-1:0] node_1220;
    wire [DATA_WIDTH-1:0] node_1221;
    wire [DATA_WIDTH-1:0] node_1222;
    wire [DATA_WIDTH-1:0] node_1223;
    wire [DATA_WIDTH-1:0] node_1224;
    wire [DATA_WIDTH-1:0] node_1225;
    wire [DATA_WIDTH-1:0] node_1226;
    wire [DATA_WIDTH-1:0] node_1227;
    wire [DATA_WIDTH-1:0] node_1228;
    wire [DATA_WIDTH-1:0] node_1229;
    wire [DATA_WIDTH-1:0] node_1230;
    wire [DATA_WIDTH-1:0] node_1231;
    wire [DATA_WIDTH-1:0] node_1232;
    wire [DATA_WIDTH-1:0] node_1233;
    wire [DATA_WIDTH-1:0] node_1234;
    wire [DATA_WIDTH-1:0] node_1235;
    wire [DATA_WIDTH-1:0] node_1236;
    wire [DATA_WIDTH-1:0] node_1237;
    wire [DATA_WIDTH-1:0] node_1238;
    wire [DATA_WIDTH-1:0] node_1239;
    wire [DATA_WIDTH-1:0] node_1240;
    wire [DATA_WIDTH-1:0] node_1241;
    wire [DATA_WIDTH-1:0] node_1242;
    wire [DATA_WIDTH-1:0] node_1243;
    wire [DATA_WIDTH-1:0] node_1244;
    wire [DATA_WIDTH-1:0] node_1245;
    wire [DATA_WIDTH-1:0] node_1246;
    wire [DATA_WIDTH-1:0] node_1247;
    wire [DATA_WIDTH-1:0] node_1248;
    wire [DATA_WIDTH-1:0] node_1249;
    wire [DATA_WIDTH-1:0] node_1250;
    wire [DATA_WIDTH-1:0] node_1251;
    wire [DATA_WIDTH-1:0] node_1252;
    wire [DATA_WIDTH-1:0] node_1253;
    wire [DATA_WIDTH-1:0] node_1254;
    wire [DATA_WIDTH-1:0] node_1255;
    wire [DATA_WIDTH-1:0] node_1256;
    wire [DATA_WIDTH-1:0] node_1257;
    wire [DATA_WIDTH-1:0] node_1258;
    wire [DATA_WIDTH-1:0] node_1259;
    wire [DATA_WIDTH-1:0] node_1260;
    wire [DATA_WIDTH-1:0] node_1261;
    wire [DATA_WIDTH-1:0] node_1262;
    wire [DATA_WIDTH-1:0] node_1263;
    wire [DATA_WIDTH-1:0] node_1264;
    wire [DATA_WIDTH-1:0] node_1265;
    wire [DATA_WIDTH-1:0] node_1266;
    wire [DATA_WIDTH-1:0] node_1267;
    wire [DATA_WIDTH-1:0] node_1268;
    wire [DATA_WIDTH-1:0] node_1269;
    wire [DATA_WIDTH-1:0] node_1270;
    wire [DATA_WIDTH-1:0] node_1271;
    wire [DATA_WIDTH-1:0] node_1272;
    wire [DATA_WIDTH-1:0] node_1273;
    wire [DATA_WIDTH-1:0] node_1274;
    wire [DATA_WIDTH-1:0] node_1275;
    wire [DATA_WIDTH-1:0] node_1276;
    wire [DATA_WIDTH-1:0] node_1277;
    wire [DATA_WIDTH-1:0] node_1278;
    wire [DATA_WIDTH-1:0] node_1279;
    wire [DATA_WIDTH-1:0] node_1280;
    wire [DATA_WIDTH-1:0] node_1281;
    wire [DATA_WIDTH-1:0] node_1282;
    wire [DATA_WIDTH-1:0] node_1283;
    wire [DATA_WIDTH-1:0] node_1284;
    wire [DATA_WIDTH-1:0] node_1285;
    wire [DATA_WIDTH-1:0] node_1286;
    wire [DATA_WIDTH-1:0] node_1287;
    wire [DATA_WIDTH-1:0] node_1288;
    wire [DATA_WIDTH-1:0] node_1289;
    wire [DATA_WIDTH-1:0] node_1290;
    wire [DATA_WIDTH-1:0] node_1291;
    wire [DATA_WIDTH-1:0] node_1292;
    wire [DATA_WIDTH-1:0] node_1293;
    wire [DATA_WIDTH-1:0] node_1294;
    wire [DATA_WIDTH-1:0] node_1295;
    wire [DATA_WIDTH-1:0] node_1296;
    wire [DATA_WIDTH-1:0] node_1297;
    wire [DATA_WIDTH-1:0] node_1298;
    wire [DATA_WIDTH-1:0] node_1299;
    wire [DATA_WIDTH-1:0] node_1300;
    wire [DATA_WIDTH-1:0] node_1301;
    wire [DATA_WIDTH-1:0] node_1302;
    wire [DATA_WIDTH-1:0] node_1303;
    wire [DATA_WIDTH-1:0] node_1304;
    wire [DATA_WIDTH-1:0] node_1305;
    wire [DATA_WIDTH-1:0] node_1306;
    wire [DATA_WIDTH-1:0] node_1307;
    wire [DATA_WIDTH-1:0] node_1308;
    wire [DATA_WIDTH-1:0] node_1309;
    wire [DATA_WIDTH-1:0] node_1310;
    wire [DATA_WIDTH-1:0] node_1311;
    wire [DATA_WIDTH-1:0] node_1312;
    wire [DATA_WIDTH-1:0] node_1313;
    wire [DATA_WIDTH-1:0] node_1314;
    wire [DATA_WIDTH-1:0] node_1315;
    wire [DATA_WIDTH-1:0] node_1316;
    wire [DATA_WIDTH-1:0] node_1317;
    wire [DATA_WIDTH-1:0] node_1318;
    wire [DATA_WIDTH-1:0] node_1319;
    wire [DATA_WIDTH-1:0] node_1320;
    wire [DATA_WIDTH-1:0] node_1321;
    wire [DATA_WIDTH-1:0] node_1322;
    wire [DATA_WIDTH-1:0] node_1323;
    wire [DATA_WIDTH-1:0] node_1324;
    wire [DATA_WIDTH-1:0] node_1325;
    wire [DATA_WIDTH-1:0] node_1326;
    wire [DATA_WIDTH-1:0] node_1327;
    wire [DATA_WIDTH-1:0] node_1328;
    wire [DATA_WIDTH-1:0] node_1329;
    wire [DATA_WIDTH-1:0] node_1330;
    wire [DATA_WIDTH-1:0] node_1331;
    wire [DATA_WIDTH-1:0] node_1332;
    wire [DATA_WIDTH-1:0] node_1333;
    wire [DATA_WIDTH-1:0] node_1334;
    wire [DATA_WIDTH-1:0] node_1335;
    wire [DATA_WIDTH-1:0] node_1336;
    wire [DATA_WIDTH-1:0] node_1337;
    wire [DATA_WIDTH-1:0] node_1338;
    wire [DATA_WIDTH-1:0] node_1339;
    wire [DATA_WIDTH-1:0] node_1340;
    wire [DATA_WIDTH-1:0] node_1341;
    wire [DATA_WIDTH-1:0] node_1342;
    wire [DATA_WIDTH-1:0] node_1343;
    wire [DATA_WIDTH-1:0] node_1344;
    wire [DATA_WIDTH-1:0] node_1345;
    wire [DATA_WIDTH-1:0] node_1346;
    wire [DATA_WIDTH-1:0] node_1347;
    wire [DATA_WIDTH-1:0] node_1348;
    wire [DATA_WIDTH-1:0] node_1349;
    wire [DATA_WIDTH-1:0] node_1350;
    wire [DATA_WIDTH-1:0] node_1351;
    wire [DATA_WIDTH-1:0] node_1352;
    wire [DATA_WIDTH-1:0] node_1353;
    wire [DATA_WIDTH-1:0] node_1354;
    wire [DATA_WIDTH-1:0] node_1355;
    wire [DATA_WIDTH-1:0] node_1356;
    wire [DATA_WIDTH-1:0] node_1357;
    wire [DATA_WIDTH-1:0] node_1358;
    wire [DATA_WIDTH-1:0] node_1359;
    wire [DATA_WIDTH-1:0] node_1360;
    wire [DATA_WIDTH-1:0] node_1361;
    wire [DATA_WIDTH-1:0] node_1362;
    wire [DATA_WIDTH-1:0] node_1363;
    wire [DATA_WIDTH-1:0] node_1364;
    wire [DATA_WIDTH-1:0] node_1365;
    wire [DATA_WIDTH-1:0] node_1366;
    wire [DATA_WIDTH-1:0] node_1367;
    wire [DATA_WIDTH-1:0] node_1368;
    wire [DATA_WIDTH-1:0] node_1369;
    wire [DATA_WIDTH-1:0] node_1370;
    wire [DATA_WIDTH-1:0] node_1371;
    wire [DATA_WIDTH-1:0] node_1372;
    wire [DATA_WIDTH-1:0] node_1373;
    wire [DATA_WIDTH-1:0] node_1374;
    wire [DATA_WIDTH-1:0] node_1375;
    wire [DATA_WIDTH-1:0] node_1376;
    wire [DATA_WIDTH-1:0] node_1377;
    wire [DATA_WIDTH-1:0] node_1378;
    wire [DATA_WIDTH-1:0] node_1379;
    wire [DATA_WIDTH-1:0] node_1380;
    wire [DATA_WIDTH-1:0] node_1381;
    wire [DATA_WIDTH-1:0] node_1382;
    wire [DATA_WIDTH-1:0] node_1383;
    wire [DATA_WIDTH-1:0] node_1384;
    wire [DATA_WIDTH-1:0] node_1385;
    wire [DATA_WIDTH-1:0] node_1386;
    wire [DATA_WIDTH-1:0] node_1387;
    wire [DATA_WIDTH-1:0] node_1388;
    wire [DATA_WIDTH-1:0] node_1389;
    wire [DATA_WIDTH-1:0] node_1390;
    wire [DATA_WIDTH-1:0] node_1391;
    wire [DATA_WIDTH-1:0] node_1392;
    wire [DATA_WIDTH-1:0] node_1393;
    wire [DATA_WIDTH-1:0] node_1394;
    wire [DATA_WIDTH-1:0] node_1395;
    wire [DATA_WIDTH-1:0] node_1396;
    wire [DATA_WIDTH-1:0] node_1397;
    wire [DATA_WIDTH-1:0] node_1398;
    wire [DATA_WIDTH-1:0] node_1399;
    wire [DATA_WIDTH-1:0] node_1400;
    wire [DATA_WIDTH-1:0] node_1401;
    wire [DATA_WIDTH-1:0] node_1402;
    wire [DATA_WIDTH-1:0] node_1403;
    wire [DATA_WIDTH-1:0] node_1404;
    wire [DATA_WIDTH-1:0] node_1405;
    wire [DATA_WIDTH-1:0] node_1406;
    wire [DATA_WIDTH-1:0] node_1407;
    wire [DATA_WIDTH-1:0] node_1408;
    wire [DATA_WIDTH-1:0] node_1409;
    wire [DATA_WIDTH-1:0] node_1410;
    wire [DATA_WIDTH-1:0] node_1411;
    wire [DATA_WIDTH-1:0] node_1412;
    wire [DATA_WIDTH-1:0] node_1413;
    wire [DATA_WIDTH-1:0] node_1414;
    wire [DATA_WIDTH-1:0] node_1415;
    wire [DATA_WIDTH-1:0] node_1416;
    wire [DATA_WIDTH-1:0] node_1417;
    wire [DATA_WIDTH-1:0] node_1418;
    wire [DATA_WIDTH-1:0] node_1419;
    wire [DATA_WIDTH-1:0] node_1420;
    wire [DATA_WIDTH-1:0] node_1421;
    wire [DATA_WIDTH-1:0] node_1422;
    wire [DATA_WIDTH-1:0] node_1423;
    wire [DATA_WIDTH-1:0] node_1424;
    wire [DATA_WIDTH-1:0] node_1425;
    wire [DATA_WIDTH-1:0] node_1426;
    wire [DATA_WIDTH-1:0] node_1427;
    wire [DATA_WIDTH-1:0] node_1428;
    wire [DATA_WIDTH-1:0] node_1429;
    wire [DATA_WIDTH-1:0] node_1430;
    wire [DATA_WIDTH-1:0] node_1431;
    wire [DATA_WIDTH-1:0] node_1432;
    wire [DATA_WIDTH-1:0] node_1433;
    wire [DATA_WIDTH-1:0] node_1434;
    wire [DATA_WIDTH-1:0] node_1435;
    wire [DATA_WIDTH-1:0] node_1436;
    wire [DATA_WIDTH-1:0] node_1437;
    wire [DATA_WIDTH-1:0] node_1438;
    wire [DATA_WIDTH-1:0] node_1439;
    wire [DATA_WIDTH-1:0] node_1440;
    wire [DATA_WIDTH-1:0] node_1441;
    wire [DATA_WIDTH-1:0] node_1442;
    wire [DATA_WIDTH-1:0] node_1443;
    wire [DATA_WIDTH-1:0] node_1444;
    wire [DATA_WIDTH-1:0] node_1445;
    wire [DATA_WIDTH-1:0] node_1446;
    wire [DATA_WIDTH-1:0] node_1447;
    wire [DATA_WIDTH-1:0] node_1448;
    wire [DATA_WIDTH-1:0] node_1449;
    wire [DATA_WIDTH-1:0] node_1450;
    wire [DATA_WIDTH-1:0] node_1451;
    wire [DATA_WIDTH-1:0] node_1452;
    wire [DATA_WIDTH-1:0] node_1453;
    wire [DATA_WIDTH-1:0] node_1454;
    wire [DATA_WIDTH-1:0] node_1455;
    wire [DATA_WIDTH-1:0] node_1456;
    wire [DATA_WIDTH-1:0] node_1457;
    wire [DATA_WIDTH-1:0] node_1458;
    wire [DATA_WIDTH-1:0] node_1459;
    wire [DATA_WIDTH-1:0] node_1460;
    wire [DATA_WIDTH-1:0] node_1461;
    wire [DATA_WIDTH-1:0] node_1462;
    wire [DATA_WIDTH-1:0] node_1463;
    wire [DATA_WIDTH-1:0] node_1464;
    wire [DATA_WIDTH-1:0] node_1465;
    wire [DATA_WIDTH-1:0] node_1466;
    wire [DATA_WIDTH-1:0] node_1467;
    wire [DATA_WIDTH-1:0] node_1468;
    wire [DATA_WIDTH-1:0] node_1469;
    wire [DATA_WIDTH-1:0] node_1470;
    wire [DATA_WIDTH-1:0] node_1471;
    wire [DATA_WIDTH-1:0] node_1472;
    wire [DATA_WIDTH-1:0] node_1473;
    wire [DATA_WIDTH-1:0] node_1474;
    wire [DATA_WIDTH-1:0] node_1475;
    wire [DATA_WIDTH-1:0] node_1476;
    wire [DATA_WIDTH-1:0] node_1477;
    wire [DATA_WIDTH-1:0] node_1478;
    wire [DATA_WIDTH-1:0] node_1479;
    wire [DATA_WIDTH-1:0] node_1480;
    wire [DATA_WIDTH-1:0] node_1481;
    wire [DATA_WIDTH-1:0] node_1482;
    wire [DATA_WIDTH-1:0] node_1483;
    wire [DATA_WIDTH-1:0] node_1484;
    wire [DATA_WIDTH-1:0] node_1485;
    wire [DATA_WIDTH-1:0] node_1486;
    wire [DATA_WIDTH-1:0] node_1487;
    wire [DATA_WIDTH-1:0] node_1488;
    wire [DATA_WIDTH-1:0] node_1489;
    wire [DATA_WIDTH-1:0] node_1490;
    wire [DATA_WIDTH-1:0] node_1491;
    wire [DATA_WIDTH-1:0] node_1492;
    wire [DATA_WIDTH-1:0] node_1493;
    wire [DATA_WIDTH-1:0] node_1494;
    wire [DATA_WIDTH-1:0] node_1495;
    wire [DATA_WIDTH-1:0] node_1496;
    wire [DATA_WIDTH-1:0] node_1497;
    wire [DATA_WIDTH-1:0] node_1498;
    wire [DATA_WIDTH-1:0] node_1499;
    wire [DATA_WIDTH-1:0] node_1500;
    wire [DATA_WIDTH-1:0] node_1501;
    wire [DATA_WIDTH-1:0] node_1502;
    wire [DATA_WIDTH-1:0] node_1503;
    wire [DATA_WIDTH-1:0] node_1504;
    wire [DATA_WIDTH-1:0] node_1505;
    wire [DATA_WIDTH-1:0] node_1506;
    wire [DATA_WIDTH-1:0] node_1507;
    wire [DATA_WIDTH-1:0] node_1508;
    wire [DATA_WIDTH-1:0] node_1509;
    wire [DATA_WIDTH-1:0] node_1510;
    wire [DATA_WIDTH-1:0] node_1511;
    wire [DATA_WIDTH-1:0] node_1512;
    wire [DATA_WIDTH-1:0] node_1513;
    wire [DATA_WIDTH-1:0] node_1514;
    wire [DATA_WIDTH-1:0] node_1515;
    wire [DATA_WIDTH-1:0] node_1516;
    wire [DATA_WIDTH-1:0] node_1517;
    wire [DATA_WIDTH-1:0] node_1518;
    wire [DATA_WIDTH-1:0] node_1519;
    wire [DATA_WIDTH-1:0] node_1520;
    wire [DATA_WIDTH-1:0] node_1521;
    wire [DATA_WIDTH-1:0] node_1522;
    wire [DATA_WIDTH-1:0] node_1523;
    wire [DATA_WIDTH-1:0] node_1524;
    wire [DATA_WIDTH-1:0] node_1525;
    wire [DATA_WIDTH-1:0] node_1526;
    wire [DATA_WIDTH-1:0] node_1527;
    wire [DATA_WIDTH-1:0] node_1528;
    wire [DATA_WIDTH-1:0] node_1529;
    wire [DATA_WIDTH-1:0] node_1530;
    wire [DATA_WIDTH-1:0] node_1531;
    wire [DATA_WIDTH-1:0] node_1532;
    wire [DATA_WIDTH-1:0] node_1533;
    wire [DATA_WIDTH-1:0] node_1534;
    wire [DATA_WIDTH-1:0] node_1535;
    wire [DATA_WIDTH-1:0] node_1536;
    wire [DATA_WIDTH-1:0] node_1537;
    wire [DATA_WIDTH-1:0] node_1538;
    wire [DATA_WIDTH-1:0] node_1539;
    wire [DATA_WIDTH-1:0] node_1540;
    wire [DATA_WIDTH-1:0] node_1541;
    wire [DATA_WIDTH-1:0] node_1542;
    wire [DATA_WIDTH-1:0] node_1543;
    wire [DATA_WIDTH-1:0] node_1544;
    wire [DATA_WIDTH-1:0] node_1545;
    wire [DATA_WIDTH-1:0] node_1546;
    wire [DATA_WIDTH-1:0] node_1547;
    wire [DATA_WIDTH-1:0] node_1548;
    wire [DATA_WIDTH-1:0] node_1549;
    wire [DATA_WIDTH-1:0] node_1550;
    wire [DATA_WIDTH-1:0] node_1551;
    wire [DATA_WIDTH-1:0] node_1552;
    wire [DATA_WIDTH-1:0] node_1553;
    wire [DATA_WIDTH-1:0] node_1554;
    wire [DATA_WIDTH-1:0] node_1555;
    wire [DATA_WIDTH-1:0] node_1556;
    wire [DATA_WIDTH-1:0] node_1557;
    wire [DATA_WIDTH-1:0] node_1558;
    wire [DATA_WIDTH-1:0] node_1559;
    wire [DATA_WIDTH-1:0] node_1560;
    wire [DATA_WIDTH-1:0] node_1561;
    wire [DATA_WIDTH-1:0] node_1562;
    wire [DATA_WIDTH-1:0] node_1563;
    wire [DATA_WIDTH-1:0] node_1564;
    wire [DATA_WIDTH-1:0] node_1565;
    wire [DATA_WIDTH-1:0] node_1566;
    wire [DATA_WIDTH-1:0] node_1567;
    wire [DATA_WIDTH-1:0] node_1568;
    wire [DATA_WIDTH-1:0] node_1569;
    wire [DATA_WIDTH-1:0] node_1570;
    wire [DATA_WIDTH-1:0] node_1571;
    wire [DATA_WIDTH-1:0] node_1572;
    wire [DATA_WIDTH-1:0] node_1573;
    wire [DATA_WIDTH-1:0] node_1574;
    wire [DATA_WIDTH-1:0] node_1575;
    wire [DATA_WIDTH-1:0] node_1576;
    wire [DATA_WIDTH-1:0] node_1577;
    wire [DATA_WIDTH-1:0] node_1578;
    wire [DATA_WIDTH-1:0] node_1579;
    wire [DATA_WIDTH-1:0] node_1580;
    wire [DATA_WIDTH-1:0] node_1581;
    wire [DATA_WIDTH-1:0] node_1582;
    wire [DATA_WIDTH-1:0] node_1583;
    wire [DATA_WIDTH-1:0] node_1584;
    wire [DATA_WIDTH-1:0] node_1585;
    wire [DATA_WIDTH-1:0] node_1586;
    wire [DATA_WIDTH-1:0] node_1587;
    wire [DATA_WIDTH-1:0] node_1588;
    wire [DATA_WIDTH-1:0] node_1589;
    wire [DATA_WIDTH-1:0] node_1590;
    wire [DATA_WIDTH-1:0] node_1591;
    wire [DATA_WIDTH-1:0] node_1592;
    wire [DATA_WIDTH-1:0] node_1593;
    wire [DATA_WIDTH-1:0] node_1594;
    wire [DATA_WIDTH-1:0] node_1595;
    wire [DATA_WIDTH-1:0] node_1596;
    wire [DATA_WIDTH-1:0] node_1597;
    wire [DATA_WIDTH-1:0] node_1598;
    wire [DATA_WIDTH-1:0] node_1599;
    wire [DATA_WIDTH-1:0] node_1600;
    wire [DATA_WIDTH-1:0] node_1601;
    wire [DATA_WIDTH-1:0] node_1602;
    wire [DATA_WIDTH-1:0] node_1603;
    wire [DATA_WIDTH-1:0] node_1604;
    wire [DATA_WIDTH-1:0] node_1605;
    wire [DATA_WIDTH-1:0] node_1606;
    wire [DATA_WIDTH-1:0] node_1607;
    wire [DATA_WIDTH-1:0] node_1608;
    wire [DATA_WIDTH-1:0] node_1609;
    wire [DATA_WIDTH-1:0] node_1610;
    wire [DATA_WIDTH-1:0] node_1611;
    wire [DATA_WIDTH-1:0] node_1612;
    wire [DATA_WIDTH-1:0] node_1613;
    wire [DATA_WIDTH-1:0] node_1614;
    wire [DATA_WIDTH-1:0] node_1615;
    wire [DATA_WIDTH-1:0] node_1616;
    wire [DATA_WIDTH-1:0] node_1617;
    wire [DATA_WIDTH-1:0] node_1618;
    wire [DATA_WIDTH-1:0] node_1619;
    wire [DATA_WIDTH-1:0] node_1620;
    wire [DATA_WIDTH-1:0] node_1621;
    wire [DATA_WIDTH-1:0] node_1622;
    wire [DATA_WIDTH-1:0] node_1623;
    wire [DATA_WIDTH-1:0] node_1624;
    wire [DATA_WIDTH-1:0] node_1625;
    wire [DATA_WIDTH-1:0] node_1626;
    wire [DATA_WIDTH-1:0] node_1627;
    wire [DATA_WIDTH-1:0] node_1628;
    wire [DATA_WIDTH-1:0] node_1629;
    wire [DATA_WIDTH-1:0] node_1630;
    wire [DATA_WIDTH-1:0] node_1631;
    wire [DATA_WIDTH-1:0] node_1632;
    wire [DATA_WIDTH-1:0] node_1633;
    wire [DATA_WIDTH-1:0] node_1634;
    wire [DATA_WIDTH-1:0] node_1635;
    wire [DATA_WIDTH-1:0] node_1636;
    wire [DATA_WIDTH-1:0] node_1637;
    wire [DATA_WIDTH-1:0] node_1638;
    wire [DATA_WIDTH-1:0] node_1639;
    wire [DATA_WIDTH-1:0] node_1640;
    wire [DATA_WIDTH-1:0] node_1641;
    wire [DATA_WIDTH-1:0] node_1642;
    wire [DATA_WIDTH-1:0] node_1643;
    wire [DATA_WIDTH-1:0] node_1644;
    wire [DATA_WIDTH-1:0] node_1645;
    wire [DATA_WIDTH-1:0] node_1646;
    wire [DATA_WIDTH-1:0] node_1647;
    wire [DATA_WIDTH-1:0] node_1648;
    wire [DATA_WIDTH-1:0] node_1649;
    wire [DATA_WIDTH-1:0] node_1650;
    wire [DATA_WIDTH-1:0] node_1651;
    wire [DATA_WIDTH-1:0] node_1652;
    wire [DATA_WIDTH-1:0] node_1653;
    wire [DATA_WIDTH-1:0] node_1654;
    wire [DATA_WIDTH-1:0] node_1655;
    wire [DATA_WIDTH-1:0] node_1656;
    wire [DATA_WIDTH-1:0] node_1657;
    wire [DATA_WIDTH-1:0] node_1658;
    wire [DATA_WIDTH-1:0] node_1659;
    wire [DATA_WIDTH-1:0] node_1660;
    wire [DATA_WIDTH-1:0] node_1661;
    wire [DATA_WIDTH-1:0] node_1662;
    wire [DATA_WIDTH-1:0] node_1663;
    wire [DATA_WIDTH-1:0] node_1664;
    wire [DATA_WIDTH-1:0] node_1665;
    wire [DATA_WIDTH-1:0] node_1666;
    wire [DATA_WIDTH-1:0] node_1667;
    wire [DATA_WIDTH-1:0] node_1668;
    wire [DATA_WIDTH-1:0] node_1669;
    wire [DATA_WIDTH-1:0] node_1670;
    wire [DATA_WIDTH-1:0] node_1671;
    wire [DATA_WIDTH-1:0] node_1672;
    wire [DATA_WIDTH-1:0] node_1673;
    wire [DATA_WIDTH-1:0] node_1674;
    wire [DATA_WIDTH-1:0] node_1675;
    wire [DATA_WIDTH-1:0] node_1676;
    wire [DATA_WIDTH-1:0] node_1677;
    wire [DATA_WIDTH-1:0] node_1678;
    wire [DATA_WIDTH-1:0] node_1679;
    wire [DATA_WIDTH-1:0] node_1680;
    wire [DATA_WIDTH-1:0] node_1681;
    wire [DATA_WIDTH-1:0] node_1682;
    wire [DATA_WIDTH-1:0] node_1683;
    wire [DATA_WIDTH-1:0] node_1684;
    wire [DATA_WIDTH-1:0] node_1685;
    wire [DATA_WIDTH-1:0] node_1686;
    wire [DATA_WIDTH-1:0] node_1687;
    wire [DATA_WIDTH-1:0] node_1688;
    wire [DATA_WIDTH-1:0] node_1689;
    wire [DATA_WIDTH-1:0] node_1690;
    wire [DATA_WIDTH-1:0] node_1691;
    wire [DATA_WIDTH-1:0] node_1692;

    // Pipeline control signals
    reg [2:0] pipeline_valid;
    reg [2:0] pipeline_counter;

    // Combinational logic for all operations
    assign node_9 = best_ask_price - best_bid_price;  // Subtraction
    assign node_11 = (32'd100 < best_bid_qty) ? 32'd1 : 32'd0;  // Less than
    assign node_12 = (32'd100 < best_ask_qty) ? 32'd1 : 32'd0;  // Less than
    assign node_14 = (node_9 == 32'd1) ? 32'd1 : 32'd0;  // Equality
    assign node_16 = (current_position == 32'd0) ? 32'd1 : 32'd0;  // Equality
    assign node_17 = (bid_queue_strong != 0) && (node_11 != 0) ? 32'd1 : 32'd0;  // Logical AND
    assign node_18 = (ask_queue_strong != 0) && (node_12 != 0) ? 32'd1 : 32'd0;  // Logical AND
    assign node_19 = (node_16 != 0) && (node_14 != 0) ? 32'd1 : 32'd0;  // Logical AND
    assign node_20 = (node_19 != 0) && (node_17 != 0) ? 32'd1 : 32'd0;  // Logical AND
    assign node_21 = (node_16 != 0) && (node_14 != 0) ? 32'd1 : 32'd0;  // Logical AND
    assign node_22 = (node_21 != 0) && (node_18 != 0) ? 32'd1 : 32'd0;  // Logical AND
    assign node_26 = (node_22 != 0) ? 32'd2 : 32'd0;  // Multiplexer
    assign node_27 = (node_20 != 0) ? 32'd1 : node_26;  // Multiplexer
    assign node_28 = (node_22 != 0) ? best_ask_price : 32'd0;  // Multiplexer
    assign node_29 = (node_20 != 0) ? best_bid_price : node_28;  // Multiplexer
    assign node_32 = (node_20 != 0) || (node_22 != 0) ? 32'd1 : 32'd0;  // Logical OR
    assign node_33 = (node_32 != 0) ? 32'd50 : 32'd0;  // Multiplexer
    assign action = node_27;  // Output assignment
    assign price = node_29;  // Output assignment
    assign quantity = node_33;  // Output assignment

    // Pipeline control
    always @(posedge ap_clk) begin
        if (!ap_rst_n) begin
            pipeline_valid <= 3'b000;
            pipeline_counter <= 3'b000;
            ap_done <= 1'b0;
        end else if (ap_start) begin
            pipeline_valid <= {pipeline_valid[1:0], 1'b1};
            pipeline_counter <= pipeline_counter + 1;
            ap_done <= pipeline_valid[2];
        end
    end

    // Control signal assignments
    assign ap_idle = ~pipeline_valid[0];
    assign ap_ready = ~pipeline_valid[0];

endmodule
